module PruebaAND(input logic a,b,
			output z); 

assign z = a & b;

endmodule
